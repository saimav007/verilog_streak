A24)
`define SIZE 40 : The value can be passed during run time also. But it can not be passed
as argument during instantiations.
parameter SIZE 40: The value can not be changed during run time. It can be passed as
argument along with module instantiations.
